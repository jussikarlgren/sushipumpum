de
den
det
de
dem
dom
också
jag
mig
mitt
min
sin
sina
mina
ju
några
vissa
även
tex
så
blir
ej
icke
inte
och
eller
på
med
deras
att
i
om
en
ett
av
vara
varit
kring
emot
från
för
före
genom
hos
ifrån
in
innan
inom
men
mellan
mot
ned
ner
nere
när
nära
omkring
ovanpå
per
på
reda
runt
sedan
som
såsom
till
tills
trots
tvärsöver
under
upp
uppför
uppåt
ur
ut
utanför
via
vid
åt
än
jag
mig
vi
oss
han
honom
hon
henne
man
sig
denna
detta
dessa
vår
vårt
våra
din
ditt
dina
deras
er
ert
era
hans
hennes
dess
vars
vad
vilken
vilket
vilka
som
sådan
sådant
sådana
samma
någon
något
några
ingen
bara
själv
är
varit
ha
har
hade
haft
ska
skall
skulle
finnas
finns
fann
funnit
bör
borde
kunna
kan
kunde
kunnat
ville
velat
där
här
dit
hit
då
nu
sedan
tillbaka
var
någorlunda
