att	3340
det	3155
och	3107
är	2623
i	2492
som	2474
vi	2098
för	2026
en	1835
på	1617
inte	1496
har	1485
om	1220
de	1202
till	1167
den	1160
av	1133
med	1092
ett	1015
jag	887
ska	844
men	818
så	768
kan	611
vill	525
man	511
sig	504
när	489
där	465
alla	445
här	437
måste	430
var	421
–	420
vara	411
nu	403
också	382
eller	363
kommer	340
hur	327
från	324
finns	318
oss	318
många	301
år	299
får	294
få	294
då	292
än	285
andra	281
mer	265
vad	264
göra	236
utan	234
bara	226
skulle	222
ta	219
detta	216
blir	215
vår	214
ha	212
han	205
upp	204
ut	203
fler	201
över	199
mycket	199
se	197
efter	197
under	194
går	193
idag	192
behöver	191
mot	191
ser	190
allt	190
sin	187
gör	182
bli	182
ni	182
nya	176
mig	174
kunna	165
därför	163
bättre	161
våra	160
in	157
land	154
sedan	151
ju	151
säger	145
hade	145
vårt	145
hon	144
